module
endmodule
