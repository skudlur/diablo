/*
*   Package for diablo
*/

`define ALU_ADD 	7'b000_0000
`define ALU_SUB 	7'b000_0001
`define ALU_AND 	7'b000_0010
`define ALU_OR 		7'b000_0011
`define ALU_XOR 	7'b000_0100

`define ALU_SLL 	7'b000_0101
`define ALU_SRL 	7'b000_0110
`define ALU_SRA 	7'b000_0111

`define ALU_SLT 	7'b000_1000
`define ALU_SLTU 	7'b000_1001
